--*************************************************************
--* This file is automatically generated test bench template  *
--* By ACTIVE-VHDL    <TBgen v1.10>. Copyright (C) ALDEC Inc. *
--*                                                           *
--* This file was generated on:           12:06 AM, 2/22/2011 *
--* Tested entity name:                               shapipe *
--* File name contains tested entity:       .\src\shapipe.vhd *
--*************************************************************

library ieee;
use work.shatypes.all;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity shapipe_tb is
end shapipe_tb;

architecture TB_ARCHITECTURE of shapipe_tb is
	-- Component declaration of the tested unit
	component shapipe
	port(
		clk : in std_logic;
		message : in word_vector(15 downto 0);
		hash : out word_vector(7 downto 0) );
end component;

	-- Stimulus signals - signals mapped to the input and inout ports of tested entity
	signal clk : std_logic;
	signal message : word_vector(15 downto 0);
	-- Observed signals - signals mapped to the output ports of tested entity
	signal hash : word_vector(7 downto 0);

	-- Add your code here ...
	signal END_SIM : BOOLEAN := FALSE;

begin

	-- Unit Under Test port map
	UUT : shapipe
		port map
			(clk => clk,
			message => message,
			hash => hash );

	-- Add your stimulus here ...
	
	stimuli: process
	begin
		-- run for a few clocks
		wait for 20ns;
		
		message(15 downto 0) <=  (x"00000000", x"00000000", x"00000000", x"00000000",
					x"00000000", x"00000000", x"00000000", x"00000000",
					x"00000000", x"00000000", x"00000000", x"00000000",
					x"00000000", x"00000000", x"00000000", x"00000000");
		wait for 660ns;
		
		END_SIM <= TRUE;
		wait;
	end process;
	
	-- generate 10ns clock
	clock: process
	begin
		if END_SIM = FALSE then
			clk <= '1';
			wait for 5 ns;
		else
			wait;
		end if;
		
		if END_SIM = FALSE then
			clk <= '0';
			wait for 5 ns;
		else
			wait;
		end if;
	end process;

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_shapipe of shapipe_tb is
	for TB_ARCHITECTURE
		for UUT : shapipe
			use entity work.shapipe(rtl);
		end for;
	end for;
end TESTBENCH_FOR_shapipe;

